* 
* ******************************************************************************
* *                                                                            *
* *                   Copyright (C) 2004-2010, Nangate Inc.                    *
* *                           All rights reserved.                             *
* *                                                                            *
* * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
* *                                                                            *
* * All trademarks, logos, software marks, and trade names (collectively the   *
* * "Marks") in this program are proprietary to Nangate or other respective    *
* * owners that have granted Nangate the right and license to use such Marks.  *
* * You are not permitted to use the Marks without the prior written consent   *
* * of Nangate or such third party that may own the Marks.                     *
* *                                                                            *
* * This file has been provided pursuant to a License Agreement containing     *
* * restrictions on its use. This file contains valuable trade secrets and     *
* * proprietary information of Nangate Inc., and is protected by U.S. and      *
* * international laws and/or treaties.                                        *
* *                                                                            *
* * The copyright notice(s) in this file does not indicate actual or intended  *
* * publication of this file.                                                  *
* *                                                                            *
* *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
* *                                                                            *
* ******************************************************************************
* 
* 
* Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
* Local time is now Fri, 3 Dec 2010, 19:32:12.
* Main process id is 27821.
*
********************************************************************************
*                                                                              *
* Cellname:   AND2_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:24:02 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 * A2)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 VSS A2 net_0 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND2_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:23:31 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND2_X2 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 * A2)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VSS A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND2_X4.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:23:29 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND2_X4 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 * A2)
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0_m2__m1 VSS A2 net_0__m0_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_x2__m0 VDD A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_x2__m1 ZN_neg A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_0 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND3_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:18:35 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 * A2) * A3)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 net_1 A2 net_0 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 VSS A3 net_1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND3_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:18:26 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND3_X2 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 * A2) * A3)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_1 A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 VSS A3 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND3_X4.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:18:25 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND3_X4 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 * A2) * A3)
M_i_4__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0_x2__m0 ZN_neg A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0_x2__m0 ZN_neg A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0_x2__m1 VDD A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0_x2__m1 VDD A3 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_3 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND4_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:13:41 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND4_X1 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=(((A1 * A2) * A3) * A4)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 net_1 A2 net_0 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 net_2 A3 net_1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_5 VSS A4 net_2 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND4_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:13:36 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND4_X2 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=(((A1 * A2) * A3) * A4)
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_1 A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_2 A3 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VSS A4 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND4_X4.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:13:34 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AND4_X4 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=(((A1 * A2) * A3) * A4)
M_i_5__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 x1 A1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 net_0__m1 A1 x1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m1 VSS A4 net_2__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN x1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS x1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 ZN x1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS x1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_9__m0 x1 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m0 VDD A3 x1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0 x1 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 VDD A1 x1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 x1 A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 VDD A2 x1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m1 x1 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m1 VDD A4 x1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN x1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD x1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 ZN x1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD x1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ANTENNA_X1.                                                      *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:30:15 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT ANTENNA_X1 A VDD VSS 
*.PININFO A:I VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI211_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:12:12 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI211_X1 A B C1 C2 ZN VDD VSS 
*.PININFO A:I B:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 * C2) + B) + A)
M_i_1 net_0 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN C1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS B ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 ZN C2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 net_1 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_2 B net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 VDD A net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI211_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:12:11 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI211_X2 A B C1 C2 ZN VDD VSS 
*.PININFO A:I B:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 * C2) + B) + A)
M_i_2__m0 ZN B VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 VSS B ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6__m0 net_2__m0_0 B net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0 VDD A net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 net_2__m1 A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 net_1 B net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 ZN C2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 net_1 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 ZN C1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 net_1 C2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI211_X4.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:12:03 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI211_X4 A B C1 C2 ZN VDD VSS 
*.PININFO A:I B:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(!(!(((C1 * C2) + B) + A)))
M_i_0 net_0 C1 ZN_3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 ZN_3 B VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VSS A ZN_3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_8_0 ZN_4 ZN_3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_8_1 VSS ZN_3 ZN_4 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_0 ZN ZN_4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_1 VSS ZN_4 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_2 ZN ZN_4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_3 VSS ZN_4 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN_3 C1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 net_1 C2 ZN_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_2 B net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 VDD A net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9_0 ZN_4 ZN_3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9_1 VDD ZN_3 ZN_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_0 ZN ZN_4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_1 VDD ZN_4 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_2 ZN ZN_4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_3 VDD ZN_4 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI21_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:18:00 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI21_X1 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A + (B1 * B2))
M_i_1 net_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN B2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 net_1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI21_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:17:40 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI21_X2 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A + (B1 * B2))
M_i_2_0_x2_1 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_0_x2_0 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_m2__m1 net_0__m0_0__m1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_m2__m1 ZN B1 net_0__m0_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_m2__m0 net_0__m0_0__m0_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_m2__m0 VSS B2 net_0__m0_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5_0_x2_0 VDD A net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_0_x2_1 net_1 A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_x2__m0 ZN B2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_x2__m1 net_1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_x2__m0 ZN B1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_x2__m1 net_1 B2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI21_X4.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:17:48 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI21_X4 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A + (B1 * B2))
M_i_2_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_2 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_3 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN B1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 VSS B2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m2 net_0__m2 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m2 ZN B1 net_0__m2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m3 net_0__m3 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m3 VSS B2 net_0__m3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5_0 VDD A net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_1 net_1 A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_2 VDD A net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_3 net_1 A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 ZN B2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0 net_1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m1 ZN B1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 net_1 B2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m2 ZN B2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m2 net_1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m3 ZN B1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m3 net_1 B2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI221_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:07:32 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 * C2) + A) + (B1 * B2))
M_i_4 net_1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 ZN B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN C1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_9 VDD B2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 net_3 B1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 net_2 A net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 ZN C2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 net_2 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI221_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:07:38 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 * C2) + A) + (B1 * B2))
M_i_2_1 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m1 net_1__m1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 ZN B1 net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_0 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7_1 net_3 A net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m1 VDD B1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m0 net_3 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m1 VDD B2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m0 net_3 B1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_0 net_2 A net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 ZN C2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 net_2 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 ZN C1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 net_2 C2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI221_X4.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:07:31 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(!(!(((C1 * C2) + A) + (B1 * B2))))
M_i_0 net_0 C1 ZN_4 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 ZN_4 A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_1 B1 ZN_4 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 VSS B2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 ZN_4 C1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_2 C2 ZN_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 net_3 A net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 VDD B1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 VDD B2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x4_0 ZN ZN_5 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x4_1 VDD ZN_5 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x4_2 ZN ZN_5 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x4_3 VDD ZN_5 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI222_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:06:07 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + (C1 * C2))
M_i_5 net_2 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN C1 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_1 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VSS B2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_11 net_4 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10 VDD C1 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 net_4 B1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 net_3 B2 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 ZN A2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_3 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI222_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:06:14 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + (C1 * C2))
M_i_5__m1 net_2__m1 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m1 ZN C1 net_2__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m0 net_2__m0_0 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m0 VSS C2 net_2__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_1__m1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 ZN B1 net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN A1 net_0__m0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_11__m0 VDD C2 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10__m0 net_4 C1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10__m1 VDD C1 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11__m1 net_4 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m1 net_3 B2 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m0 net_4 B1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m1 net_3 B1 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m0 net_4 B2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 ZN A1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 net_3 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 ZN A2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0 net_3 A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI222_X4.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:05:54 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(!(!(((A1 * A2) + (B1 * B2)) + (C1 * C2))))
M_i_0 net_0 A1 ZN_5 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 ZN_5 B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_2 C1 ZN_5 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VSS C2 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x2_0 ZN_6 ZN_5 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x2_1 VSS ZN_5 ZN_6 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_1 VSS ZN_6 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_2 ZN ZN_6 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6 ZN_5 A1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 net_3 A2 ZN_5 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 net_4 B2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 net_3 B1 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10 net_4 C1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11 VDD C2 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_1 ZN ZN_6 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_0 VDD ZN_6 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI22_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:12:48 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI22_X1 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) + (B1 * B2))
M_i_3 net_1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 ZN B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 VDD B2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_2 B1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 ZN A1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 net_2 A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI22_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:12:55 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI22_X2 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) + (B1 * B2))
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI22_X4.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:13:02 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT AOI22_X4 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) + (B1 * B2))
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m2 net_1__m2 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m2 ZN B1 net_1__m2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m3 net_1__m3 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m3 VSS B2 net_1__m3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m2 net_0__m2 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m3 VSS A2 net_0__m3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m2 VDD B2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m2 net_2 B1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m3 VDD B1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m3 net_2 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m2 ZN A2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m2 net_2 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m3 ZN A1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m3 net_2 A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:29:49 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X1 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2 VSS A Z_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VDD A Z_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X16.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:29:14 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X16 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2_0 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_2 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_3 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_4 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_5 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_6 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_7 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_0 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_1 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_2 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_3 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_4 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_5 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_6 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_7 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:29:48 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X2 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x2_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x2_1 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x2_0 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x2_1 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X32.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:31:57 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X32 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2_0 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_2 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_3 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_4 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_5 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_6 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_7 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_8 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_9 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_10 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_11 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_12 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_13 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_14 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_15 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_16 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_17 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_18 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_19 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_20 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_21 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_22 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_23 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_24 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_25 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_26 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_27 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_28 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_29 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_30 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_31 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_0 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_1 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_2 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_3 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_4 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_5 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_6 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_7 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_8 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_9 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_10 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_11 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_12 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_13 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_14 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_15 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_16 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_17 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_18 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_19 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_20 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_21 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_22 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_23 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_24 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_25 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_26 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_27 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_28 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_29 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_30 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_31 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X4.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:29:14 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X4 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2_0 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_0 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_1 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X8.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:28:36 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X8 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2_0 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_2 Z_neg A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_3 VSS A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_0 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_1 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_2 Z_neg A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_3 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:27:46 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X1 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2 VSS A Z_neg VSS NMOS_VTL W=0.095000U L=0.050000U
M_i_0 Z Z_neg VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_3 VDD A Z_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:27:41 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X2 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2 VSS A Z_neg VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_3 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X3.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:27:23 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X3 A Z VDD VSS 
*.PININFO A:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_2_1 VSS A Z_neg VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_3_1 VDD A Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATETST_X1.                                                   *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:04:40 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATETST_X1 CK E SE GCK VDD VSS 
*.PININFO CK:I E:I SE:I GCK:O VDD:P VSS:G 
M_i_0 net_000 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 VSS E net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_001 net_000 VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_27 VSS net_004 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_39 VSS net_006 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_33 net_004 net_002 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_46 net_006 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_52 net_008 CK net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_57 VSS net_002 net_008 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_63 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_69 net_009 SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_74 VDD E net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_80 net_010 net_000 VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_95 VDD net_004 net_011 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_107 VDD net_006 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_101 net_004 net_002 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_114 net_006 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_120 net_007 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_127 VDD net_002 net_007 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_133 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATETST_X2.                                                   *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:03:58 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATETST_X2 CK E SE GCK VDD VSS 
*.PININFO CK:I E:I SE:I GCK:O VDD:P VSS:G 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 VSS E net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 net_000 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_001 net_000 VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_27 VSS net_004 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_33 net_004 net_002 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_57 VSS net_002 net_008 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_52 net_008 CK net_007 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_63 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_46 net_006 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_107 VDD net_006 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_74 VDD E net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_69 net_009 SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_80 net_010 net_000 VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_95 VDD net_004 net_011 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_101 net_004 net_002 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_127 VDD net_002 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_120 net_007 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_114 net_006 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATETST_X4.                                                   *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:03:50 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATETST_X4 CK E SE GCK VDD VSS 
*.PININFO CK:I E:I SE:I GCK:O VDD:P VSS:G 
M_i_0 net_000 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 VSS E net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_39 VSS net_006 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_001 net_000 VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_27 VSS net_004 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_33 net_004 net_002 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_46 net_006 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_52 net_008 CK VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_52_76 net_008b CK VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_63 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_69 net_009 SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_74 VDD E net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_107 VDD net_006 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_80 net_010 net_000 VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_95 VDD net_004 net_011 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_101 net_004 net_002 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_114 net_006 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_120 net_007 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_127 VDD net_002 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_120_72 net_007 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATETST_X8.                                                   *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:04:07 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATETST_X8 CK E SE GCK VDD VSS 
*.PININFO CK:I E:I SE:I GCK:O VDD:P VSS:G 
M_i_0 net_000 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 VSS E net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_39 VSS net_006 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_001 net_000 VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_27 VSS net_004 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_33_93 net_004 net_002 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_33 net_004 net_002 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_46 net_006 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_52 net_008 CK VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_52_76 net_008b CK VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_52_150 net_008c CK VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_57_123 net_007 net_002 net_008c VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_57_77_169 net_007 net_002 net_008d VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_52_76_137 net_008d CK VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_63 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_12 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_13_55 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_15_27 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_63_13_29_4 GCK net_007 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_69 net_009 SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_74 VDD E net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_107 VDD net_006 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_80 net_010 net_000 VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_95 VDD net_004 net_011 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_101_94 net_004 net_002 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_101 net_004 net_002 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_114 net_006 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_120 net_007 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_127 VDD net_002 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_120_72 net_007 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_120_163 net_007 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_127_158 VDD net_002 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_127_69_164 VDD net_002 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_120_72_145 net_007 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_38 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_10_20 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_11_14 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_133_10_28_7 GCK net_007 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATE_X1.                                                      *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:03:07 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATE_X1 CK E GCK VDD VSS 
*.PININFO CK:I E:I GCK:O VDD:P VSS:G 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_21 VSS E net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_27 net_004 net_005 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_33 VSS CK net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 VSS net_000 net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_007 CK net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_51 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_57 VDD net_002 net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_64 net_008 net_000 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_78 VDD E net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_84 net_004 net_005 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_90 VDD CK net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_103 VDD net_000 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_97 net_006 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_109 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATE_X2.                                                      *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:02:42 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATE_X2 CK E GCK VDD VSS 
*.PININFO CK:I E:I GCK:O VDD:P VSS:G 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_21 VSS E net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_27 net_004 net_005 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_33 VSS CK net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_007 CK net_006 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_45 VSS net_000 net_007 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_51 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_57 VDD net_002 net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_78 VDD E net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_64 net_008 net_000 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_84 net_004 net_005 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_90 VDD CK net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_97 net_006 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_103 VDD net_000 net_006 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATE_X4.                                                      *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:02:49 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATE_X4 CK E GCK VDD VSS 
*.PININFO CK:I E:I GCK:O VDD:P VSS:G 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_21 VSS E net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_27 net_004 net_005 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_33 VSS CK net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 VSS net_000 net_007b VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_40 net_007b CK net_006 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_51 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_57 VDD net_002 net_000 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_78 VDD E net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_64 net_008 net_000 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_84 net_004 net_005 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_90 VDD CK net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_103 VDD net_000 net_006 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_97 net_006 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_97_71 net_006 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKGATE_X8.                                                      *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:02:20 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT CLKGATE_X8 CK E GCK VDD VSS 
*.PININFO CK:I E:I GCK:O VDD:P VSS:G 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_21 VSS E net_003 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_0 VSS net_002 net_000 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_174 VSS net_002 net_000 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_33 VSS CK net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 VSS net_000 net_007b VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_40 net_007b CK net_006 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_45_63 VSS net_000 net_007c VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_40_71 net_007c CK net_006 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_40_75_82 net_007d CK net_006 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_45_66_78 VSS net_000 net_007d VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_51 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_40 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_7_58 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_10_28 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_51_7_25_30 GCK net_006 VSS VSS NMOS_VTL W=0.195000U L=0.050000U
M_i_84 net_004 net_005 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_78 VDD E net_009 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_64 net_008 net_000 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_57 VDD net_002 net_000 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_57_165 VDD net_002 net_000 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_90 VDD CK net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_103 VDD net_000 net_006 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_97 net_006 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_97_71 net_006 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_103_72 VDD net_000 net_006 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_97_99 net_006 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_97_71_87 net_006 CK VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_103_74_97 VDD net_000 net_006 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_53 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_4_22 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_24_52 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_109_4_19_36 GCK net_006 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRS_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:01:54 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFFRS_X1 D RN SN CK Q QN VDD VSS 
*.PININFO D:I RN:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_MN81 QN z99 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL W=0.210000U L=0.050000U
M_transistor_1 nn99 SN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN51 VSS z41 nn5 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN52 nn5 RN z56 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN63 VSS SN nn62 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN62 nn62 z56 nn61 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN41 z41 ck_i nn4 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN42 nn4 z37 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MP91_1 nn2 SN z51 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN33 VSS RN nn32 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN32 nn32 z51 nn31 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN31 nn31 ck_i z37 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN12 nn1 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN91 ckn_i CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MP81_0 QN z99 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP81_1 VDD z56 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_transistor_2 VDD z56 z99 VDD PMOS_VTL W=0.315000U L=0.050000U
M_transistor_3 z99 SN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP51 z56 z41 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP52 VDD RN z56 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP63 VDD SN np61 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP61 VDD z56 np61 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP62 np61 ck_i z41 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP41 np4 ckn_i z41 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP42 VDD z37 np4 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP21 VDD z37 z51 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP22 z51 SN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP33 VDD RN np32 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP31 VDD z51 np32 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP34 np32 ckn_i z37 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP12 np1 ck_i z37 VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP11 VDD D np1 VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP91 ckn_i CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRS_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:01:53 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFFRS_X2 D RN SN CK Q QN VDD VSS 
*.PININFO D:I RN:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_MN81_53 QN z99 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN81 QN z99 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN91_0_0_58 VSS z56 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL W=0.310000U L=0.050000U
M_transistor_1 nn99 SN VSS VSS NMOS_VTL W=0.310000U L=0.050000U
M_MN51 VSS RN nn5 VSS NMOS_VTL W=0.310000U L=0.050000U
M_MN52 nn5 z41 z56 VSS NMOS_VTL W=0.310000U L=0.050000U
M_MN63 VSS SN nn62 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN62 nn62 z56 nn61 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN41 z41 ck_i nn4 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN42 nn4 z37 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MP91_1 nn2 SN z51 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN33 VSS RN nn32 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN32 nn32 z51 nn31 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN31 nn31 ck_i z37 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN12 nn1 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN91 ckn_i CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MP81_0_51 QN z99 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP81_0 QN z99 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP81_1 VDD z56 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP81_1_55 VDD z56 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_transistor_2 VDD z56 z99 VDD PMOS_VTL W=0.485000U L=0.050000U
M_transistor_3 z99 SN VDD VDD PMOS_VTL W=0.485000U L=0.050000U
M_MP52 VDD RN z56 VDD PMOS_VTL W=0.485000U L=0.050000U
M_MP51 z56 z41 VDD VDD PMOS_VTL W=0.485000U L=0.050000U
M_MP63 VDD SN np61 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP61 VDD z56 np61 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP62 np61 ck_i z41 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP41 np4 ckn_i z41 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP42 VDD z37 np4 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP21 VDD z37 z51 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP22 z51 SN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP33 VDD RN np32 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP31 VDD z51 np32 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP34 np32 ckn_i z37 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP12 np1 ck_i z37 VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP11 VDD D np1 VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP91 ckn_i CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFR_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:01:01 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFFR_X1 D RN CK Q QN VDD VSS 
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_0 VSS CK net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_32 VSS RN net_005 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_38 VSS net_003 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 net_007 net_003 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_59 VSS net_011 net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_65 net_010 RN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_76 VSS net_008 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_83 Q net_011 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_89 VDD CK net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_96 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_103 net_012 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_119 VDD net_006 net_013 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_125 net_013 RN VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_136 VDD net_003 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_143 net_015 net_003 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_159 VDD net_011 net_016 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_165 net_011 RN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_172 VDD net_008 net_011 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_180 VDD net_008 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_187 Q net_011 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFR_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:00:47 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFFR_X2 D RN CK Q QN VDD VSS 
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_0 VSS CK net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_32 VSS RN net_005 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_38 VSS net_003 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 net_007 net_003 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_59 VSS net_011 net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_65 net_010 RN VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_76_4 VSS net_008 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_76 VSS net_008 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_83 Q net_011 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_83_49 Q net_011 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_89 VDD CK net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_96 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_103 net_012 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_119 VDD net_006 net_013 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_125 net_013 RN VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_136 VDD net_003 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_143 net_015 net_003 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_159 VDD net_011 net_016 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_165 net_011 RN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_172 VDD net_008 net_011 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_180_3 VDD net_008 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_180 VDD net_008 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_187 Q net_011 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_187_39 Q net_011 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFS_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:00:41 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFFS_X1 D SN CK Q QN VDD VSS 
*.PININFO D:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_15 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_30 VSS net_006 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_36 net_005 SN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 VSS CK net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_73 VSS net_003 net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_53 net_008 SN VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_46 VSS net_010 net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_86 QN net_010 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_79 VSS net_007 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_99 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_106 net_012 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_122 VDD net_006 net_013 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_128 net_006 SN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_134 VDD net_003 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_92 VDD CK net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_171 net_016 net_003 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_165 VDD net_007 net_015 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_149 net_015 SN VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_142 VDD net_010 net_007 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_189 QN net_010 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_182 VDD net_007 Q VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFS_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:00:00 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFFS_X2 D SN CK Q QN VDD VSS 
*.PININFO D:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_15 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_30 VSS net_006 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_36 net_005 SN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 VSS CK net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_73 VSS net_003 net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_53 net_008 SN VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_79_29 VSS net_007 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_79 VSS net_007 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_86 QN net_010 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_86_15 QN net_010 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_46 VSS net_010 net_007 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_99 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_106 net_012 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_122 VDD net_006 net_013 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_128 net_006 SN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_134 VDD net_003 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_92 VDD CK net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_171 net_016 net_003 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_165 VDD net_007 net_015 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_149 net_015 SN VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_182_20 VDD net_007 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_182 VDD net_007 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_189 QN net_010 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_189_10 QN net_010 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_142 VDD net_010 net_007 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFF_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:59:45 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFF_X1 D CK Q QN VDD VSS 
*.PININFO D:I CK:I Q:O QN:O VDD:P VSS:G 
M_MN2 ci cni VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN6 VSS z4 z6 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN7 z3 ci z6 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN4 z2 cni z3 VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN3 z2 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN5 z4 z3 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN1 VSS CK cni VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN8 z12 z3 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN9 z9 ci z12 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN12 z9 cni z8 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN11 z8 z10 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN10 VSS z9 z10 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN14 QN z9 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN13 VSS z10 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_MP2 ci cni VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP6 VDD z4 z1 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP7 z1 cni z3 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP4 z3 ci z5 VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP3 z5 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP5 z4 z3 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP1 VDD CK cni VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP8 z7 z3 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP9 z9 cni z7 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP12 z9 ci z11 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP11 z11 z10 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP10 VDD z9 z10 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP14 QN z9 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP13 VDD z10 Q VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFF_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:59:42 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DFF_X2 D CK Q QN VDD VSS 
*.PININFO D:I CK:I Q:O QN:O VDD:P VSS:G 
M_MN2 ci cni VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN6 VSS z4 z6 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN7 z3 ci z6 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN4 z2 cni z3 VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN3 z2 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_MN5 z4 z3 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN1 VSS CK cni VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN8 z12 z3 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN9 z9 ci z12 VSS NMOS_VTL W=0.210000U L=0.050000U
M_MN12 z9 cni z8 VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN11 z8 z10 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_MN10 VSS z9 z10 VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN14_8 QN z9 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN14 QN z9 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN13 VSS z10 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_MN13_38 VSS z10 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_MP2 ci cni VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP6 VDD z4 z1 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP7 z1 cni z3 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP4 z3 ci z5 VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP3 z5 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_MP5 z4 z3 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP1 VDD CK cni VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP8 z7 z3 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP9 z9 cni z7 VDD PMOS_VTL W=0.315000U L=0.050000U
M_MP12 z9 ci z11 VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP11 z11 z10 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_MP10 VDD z9 z10 VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP14_5 QN z9 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP14 QN z9 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP13 VDD z10 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_MP13_26 VDD z10 Q VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLH_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:59:00 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DLH_X1 D G Q VDD VSS 
*.PININFO D:I G:I Q:O VDD:P VSS:G 
M_i_0 VSS G net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_41_11 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_28 VSS net_005 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_34 VSS net_003 net_005 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_48 VDD G net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_89_4 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_55 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_61 net_006 D VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_76 VDD net_005 net_007 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_82 VDD net_003 net_005 VDD PMOS_VTL W=0.090000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLH_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:58:52 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DLH_X2 D G Q VDD VSS 
*.PININFO D:I G:I Q:O VDD:P VSS:G 
M_i_0 VSS G net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_41 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_41_11 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_28 VSS net_005 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_34 VSS net_003 net_005 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_48 VDD G net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_89 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_89_4 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_55 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_61 net_006 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_76 VDD net_005 net_007 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_82 VDD net_003 net_005 VDD PMOS_VTL W=0.090000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLL_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:58:46 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DLL_X1 D GN Q VDD VSS 
*.PININFO D:I GN:I Q:O VDD:P VSS:G 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_29 VSS net_005 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_35 VSS net_003 net_005 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_42 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_000 GN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_55 VDD net_000 net_001 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_62 net_006 D VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_79 VDD net_005 net_007 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_85 VDD net_003 net_005 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_92 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_48 net_000 GN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLL_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:58:19 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT DLL_X2 D GN Q VDD VSS 
*.PININFO D:I GN:I Q:O VDD:P VSS:G 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_29 VSS net_005 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_35 VSS net_003 net_005 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_42_3 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_42 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_000 GN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_55 VDD net_000 net_001 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_62 net_006 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_79 VDD net_005 net_007 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_85 VDD net_003 net_005 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_92_11 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_92 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_48 net_000 GN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FA_X1.                                                           *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:17:24 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT FA_X1 A B CI CO S VDD VSS 
*.PININFO A:I B:I CI:I CO:O S:O VDD:P VSS:G 
*.EQN CO=((A * B) + (CI * (A + B)));S=(CI ^ (A ^ B))
M_instance_159 CO net_001 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_instance_166 VSS B net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_170 net_000 A net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_176 net_001 CI net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_188 net_002 A VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_182 VSS B net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_227 net_006 B VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_215 VSS CI net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_221 net_006 A VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_209 net_005 net_001 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_203 net_004 CI net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_199 net_003 B net_004 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_194 VSS A net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_instance_233 S net_005 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_instance_239 CO net_001 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_instance_246 VDD B net_007 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_251 net_007 A net_001 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_257 net_001 CI net_008 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_269 net_008 A VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_263 VDD B net_008 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_309 net_011 B VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_297 VDD CI net_011 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_303 net_011 A VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_290 net_005 net_001 net_011 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_284 net_010 CI net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_280 net_009 B net_010 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_275 VDD A net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_instance_315 S net_005 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   WELLTAP_X1.                                                      *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Handwritten by Christopher Torng, clt67@cornell.edu                          *
*                                                                              *
********************************************************************************
.SUBCKT WELLTAP_X1 VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCELL_X1.                                                     *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:27:14 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT FILLCELL_X1 VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCELL_X16.                                                    *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:26:23 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT FILLCELL_X16 VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCELL_X2.                                                     *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:27:07 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT FILLCELL_X2 VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCELL_X32.                                                    *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:26:13 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT FILLCELL_X32 VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCELL_X4.                                                     *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:26:50 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT FILLCELL_X4 VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCELL_X8.                                                     *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:26:40 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT FILLCELL_X8 VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   HA_X1.                                                           *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:23:27 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT HA_X1 A B CO S VDD VSS 
*.PININFO A:I B:I CO:O S:O VDD:P VSS:G 
*.EQN CO=(A * B);S=(A ^ B)
M_i_1 net_0 B VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 S A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS x1 S VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 x1 B VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_6 VSS A x1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_12 net_3 A CO_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 VSS B net_3 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_10 CO CO_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 S B net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 net_1 A S VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD x1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 net_2 B VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_8 x1 A net_2 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_14 CO_neg A VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_15 VDD B CO_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_11 CO CO_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:25:52 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT INV_X1 A ZN VDD VSS 
*.PININFO A:I ZN:O VDD:P VSS:G 
*.EQN ZN=!A
M_i_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X16.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:25:12 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT INV_X16 A ZN VDD VSS 
*.PININFO A:I ZN:O VDD:P VSS:G 
*.EQN ZN=!A
M_i_0_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_4 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_5 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_6 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_7 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_8 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_9 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_10 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_11 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_12 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_13 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_4 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_5 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_6 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_7 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_8 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_9 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_10 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_11 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_12 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_13 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_14 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_15 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:25:46 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT INV_X2 A ZN VDD VSS 
*.PININFO A:I ZN:O VDD:P VSS:G 
*.EQN ZN=!A
M_i_0_0_x2_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x2_1 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_0_x2_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x2_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X32.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:26:38 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT INV_X32 A ZN VDD VSS 
*.PININFO A:I ZN:O VDD:P VSS:G 
*.EQN ZN=!A
M_i_0_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_4 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_5 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_6 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_7 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_8 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_9 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_10 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_11 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_12 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_13 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_16 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_17 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_18 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_19 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_20 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_21 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_22 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_23 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_24 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_25 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_26 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_27 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_28 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_29 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_30 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_31 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_4 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_5 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_6 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_7 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_8 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_9 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_10 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_11 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_12 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_13 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_14 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_15 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_16 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_17 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_18 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_19 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_20 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_21 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_22 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_23 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_24 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_25 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_26 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_27 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_28 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_29 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_30 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_31 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X4.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:25:21 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT INV_X4 A ZN VDD VSS 
*.PININFO A:I ZN:O VDD:P VSS:G 
*.EQN ZN=!A
M_i_0_0_x4_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_1 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_2 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_3 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_0_x4_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_2 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_3 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X8.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:24:46 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT INV_X8 A ZN VDD VSS 
*.PININFO A:I ZN:O VDD:P VSS:G 
*.EQN ZN=!A
M_i_0_0_x8_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x8_1 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x8_2 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x8_3 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x8_4 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x8_5 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x8_6 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x8_7 VSS A ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_0_x8_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x8_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x8_2 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x8_3 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x8_4 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x8_5 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x8_6 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x8_7 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LOGIC0_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:24:00 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT LOGIC0_X1 Z VDD VSS 
*.PININFO Z:O VDD:P VSS:G 
M_n_tran_1 VSS A Z VSS NMOS_VTL W=0.090000U L=0.050000U
M_transistor_0 VDD A A VDD PMOS_VTL W=0.090000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LOGIC1_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:23:59 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT LOGIC1_X1 Z VDD VSS 
*.PININFO Z:O VDD:P VSS:G 
M_n_tran_1 VSS A A VSS NMOS_VTL W=0.090000U L=0.050000U
M_p_tran_2 VDD A Z VDD PMOS_VTL W=0.135000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX2_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:17:01 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT MUX2_X1 A B S Z VDD VSS 
*.PININFO A:I B:I S:I Z:O VDD:P VSS:G 
*.EQN Z=((S * B) + (A * !S))
M_i_10 VSS S x1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 net_1 A VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_5 Z_neg x1 net_1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_2 Z_neg S net_0 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 net_0 B VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_11 VDD S x1 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_8 VDD A net_2 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_6 net_2 S Z_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_9 net_3 x1 Z_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 VDD B net_3 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX2_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:16:57 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT MUX2_X2 A B S Z VDD VSS 
*.PININFO A:I B:I S:I Z:O VDD:P VSS:G 
*.EQN Z=((S * B) + (A * !S))
M_i_4 net_1 A Z_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VSS x1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_0 B VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 Z_neg S net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10 VSS S x1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_8 VDD A net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 net_2 x1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 Z_neg B net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_2 S Z_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 VDD Z_neg Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 Z Z_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11 VDD S x1 VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND2_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:22:54 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 * A2)
M_i_1 net_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND2_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:22:47 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND2_X2 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 * A2)
M_i_1__m0_m2__m0 net_0__m0__m0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_m2__m0 ZN A1 net_0__m0__m0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_m2__m1 net_0__m0__m1 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_m2__m1 VSS A2 net_0__m0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0_x2__m0 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_x2__m0 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_x2__m1 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_x2__m1 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND2_X4.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:22:44 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND2_X4 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 * A2)
M_i_1_0 VSS A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_1 net_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_2 VSS A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_3 net_0 A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_0 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_1 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_2 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_3 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2_0 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2_1 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2_2 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2_3 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND3_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:16:24 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) * A3)
M_i_2 net_1 A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 ZN A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND3_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:16:17 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND3_X2 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) * A3)
M_i_2__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_m2__m0 ZN A1 net_0__m0_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_m2__m1 net_0__m0_0__m1 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m0_x2__m0 ZN A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_x2__m0 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_x2__m0 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_x2__m1 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_x2__m1 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0_x2__m1 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND3_X4.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:16:27 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND3_X4 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 * A2) * A3)
M_i_2__m0 net_1__m0_0 A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 VSS A3 net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m2 net_1__m2 A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m2 net_0__m2 A2 net_1__m2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m3 net_1__m3 A2 net_0__m3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m3 VSS A3 net_1__m3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m0 ZN A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m1 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m2 ZN A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m2 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m2 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m3 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m3 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m3 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND4_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:11:28 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND4_X1 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 * A2) * A3) * A4)
M_i_3 net_2 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_1 A3 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 ZN A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND4_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:11:18 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND4_X2 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 * A2) * A3) * A4)
M_i_3__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 VSS A4 net_2__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0 ZN A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 ZN A1 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 VDD A2 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 ZN A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 VDD A4 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND4_X4.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:11:34 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NAND4_X4 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 * A2) * A3) * A4)
M_i_0_187 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_85 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_34 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_177 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_24 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_75 net_0 A2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_196 net_1 A3 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_94 net_1 A3 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_43 net_1 A3 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_1 A3 net_2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_170 net_2 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_68 net_2 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_17 net_2 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_2 A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4_168 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_66 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_15 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 VDD A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_189 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_36 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_87 ZN A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6_202 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6_100 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6_49 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 VDD A3 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_154 ZN A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_52 ZN A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_1 ZN A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 ZN A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR2_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:22:22 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 + A2)
M_i_1 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_0 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR2_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:22:11 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR2_X2 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 + A2)
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR2_X4.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:22:01 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR2_X4 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A1 + A2)
M_i_1__m0_x2__m0_16 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_x2__m0_35 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_x2__m1_57 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_x2__m1_23 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0_m2__m0_38 net_0__m0__m3 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_m2__m0_52 ZN A1 net_0__m0__m3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_m2__m1_45 net_0__m0__m2 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_m2__m1_58 VDD A2 net_0__m0__m2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR3_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:15:39 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) + A3)
M_i_2 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 net_1 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR3_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:15:33 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR3_X2 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) + A3)
M_i_2_0_x2__m0 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_1_x2__m0 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x2__m0 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x2__m1 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_1_x2__m1 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_0_x2__m1 VSS A3 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5_1_m2__m0 net_1_0__m0_0 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_0_m2__m0 net_0_0__m0_0 A2 net_1_0__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_1_m2__m0 ZN A1 net_0_0__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_1_m2__m1 net_0_0__m1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_0_m2__m1 net_1_0__m1 A2 net_0_0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_1_m2__m1 VDD A3 net_1_0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR3_X4.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:15:48 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR3_X4 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) + A3)
M_i_0_28 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_19 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_10 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_31 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_40 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_49 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_58 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_67 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_85 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_24 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_15 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3_6 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_34 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_43 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_52 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 net_1 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_56 net_1 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_65 net_1 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_83 net_1 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR4_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:10:34 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR4_X1 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) + A4)
M_i_3 ZN A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS A3 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 net_2 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_1 A3 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR4_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:10:31 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR4_X2 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) + A4)
M_i_3__m0 ZN A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 VSS A3 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 VSS A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 ZN A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 VSS A4 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 ZN A1 net_0__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 net_0__m1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 VDD A4 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR4_X4.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:10:50 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT NOR4_X4 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) + A4)
M_i_0_22 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_22_71 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_77 VSS A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_13 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_13_89 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1_79 ZN A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS A3 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_29 VSS A3 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_52 VSS A3 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_29_45 VSS A3 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 ZN A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_8 ZN A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_109 ZN A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3_8_108 ZN A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4_6 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_6_75 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4_68 ZN A1 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_24 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_24_95 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_88 net_0 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_1 A3 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6_34 net_1 A3 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6_56 net_1 A3 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6_34_44 net_1 A3 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 net_2 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_1 net_2 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_102 net_2 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_1_96 net_2 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI211_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:09:02 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI211_X1 A B C1 C2 ZN VDD VSS 
*.PININFO A:I B:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 + C2) * A) * B)
M_i_1 ZN C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_0 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_1 A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VSS B net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 net_2 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 ZN C1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 ZN B VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI211_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:08:59 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI211_X2 A B C1 C2 ZN VDD VSS 
*.PININFO A:I B:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 + C2) * A) * B)
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6__m0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0 VDD B ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 ZN B VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI211_X4.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:09:10 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI211_X4 A B C1 C2 ZN VDD VSS 
*.PININFO A:I B:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 + C2) * A) * B)
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m2 net_1__m2 A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m2 VSS B net_1__m2 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m3 net_1__m3 B VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m3 net_0 A net_1__m3 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m2 ZN C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m2 net_0 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m3 ZN C1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m3 net_0 C2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6__m0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0 VDD B ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 ZN B VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m2 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m2 VDD B ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m3 ZN B VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m3 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m2 net_2__m2 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m2 ZN C1 net_2__m2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m3 net_2__m3 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m3 VDD C2 net_2__m3 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI21_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:14:54 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI21_X1 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A * (B1 + B2))
M_i_1 ZN B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 VSS A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_1 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3 ZN B1 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI21_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:14:55 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI21_X2 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A * (B1 + B2))
M_i_2_0 VSS A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 net_0 A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI21_X4.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:15:03 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI21_X4 A B1 B2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A * (B1 + B2))
M_i_2_0 VSS A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 net_0 A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_2 VSS A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_3 net_0 A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m2 ZN B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m2 net_0 B1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m3 ZN B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m3 net_0 B2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_2 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5_3 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m2 net_1__m2 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m2 ZN B1 net_1__m2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_3__m3 net_1__m3 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m3 VDD B2 net_1__m3 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI221_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:06:54 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 + C2) * A) * (B1 + B2))
M_i_4 VSS B2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_1 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_0 A net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 ZN C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_0 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_9 net_3 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 ZN B1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_2 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 ZN C1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI221_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:06:53 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((C1 + C2) * A) * (B1 + B2))
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_1 net_1 A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 VSS B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m1 net_1 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m0 VSS B2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_1 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2_0 net_0 A net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 net_2__m1 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 VDD C2 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_0 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7_1 VDD A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI221_X4.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:06:43 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(!(!(((C1 + C2) * A) * (B1 + B2))))
M_i_0 ZN_4 C1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 C2 ZN_4 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_1 A net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VSS B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 VSS B2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 net_2 C1 ZN_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 VDD C2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 ZN_4 A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 net_3 B1 ZN_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 VDD B2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_3_x4_3 ZN ZN_5 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_3_x4_2 VDD ZN_5 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_3_x4_1 ZN ZN_5 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_3_x4_0 VDD ZN_5 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI222_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:05:21 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * (C1 + C2))
M_i_5 net_1 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 VSS C1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_1 B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_0 B2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 ZN A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_11 net_4 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10 ZN C1 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 net_3 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 VDD B2 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 net_2 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 ZN A1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI222_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:05:02 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * (C1 + C2))
M_i_4__m0 VSS C1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m1 net_1 C2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m0 VSS C2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m1 net_1 C1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 net_0 B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 net_1 B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_0 B2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 net_1 B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_10__m1 net_4__m1 C1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11__m1 VDD C2 net_4__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11__m0 net_4__m0_0 C2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10__m0 ZN C1 net_4__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 net_2__m0_0 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0 VDD A2 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 net_2__m1 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 ZN A1 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI222_X4.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:04:48 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(!(!(((A1 + A2) * (B1 + B2)) * (C1 + C2))))
M_i_0 ZN_5 A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 ZN_5 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_1 B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_0 B1 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_1 C1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VSS C2 net_1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_1_x2_1 ZN_6 ZN_5 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_12_1_x2_0 VSS ZN_5 ZN_6 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_2 VSS ZN_6 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_1 ZN ZN_6 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6 net_2 A1 ZN_5 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 VDD A2 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 net_3 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 ZN_5 B1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10 net_4 C1 ZN_5 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_11 VDD C2 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_0 ZN ZN_6 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_15_3_x4_1 VDD ZN_6 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI22_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:09:49 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI22_X1 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) * (B1 + B2))
M_i_3 VSS B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 net_0 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 net_2 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 ZN B1 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4 net_1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI22_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:09:44 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI22_X2 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) * (B1 + B2))
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI22_X4.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:09:56 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI22_X4 A1 A2 B1 B2 ZN VDD VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VSS:G 
*.EQN ZN=!((A1 + A2) * (B1 + B2))
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m2 VSS B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m2 net_0 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m3 VSS B1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m3 net_0 B2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m2 ZN A2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m2 net_0 A1 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0__m3 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1__m3 net_0 A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m2 net_2__m2 B2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m2 ZN B1 net_2__m2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m3 net_2__m3 B1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m3 VDD B2 net_2__m3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m2 net_1__m2 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m2 ZN A1 net_1__m2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m3 net_1__m3 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m3 VDD A2 net_1__m3 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI33_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:05:27 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OAI33_X1 A1 A2 A3 B1 B2 B3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * ((B1 + B2) + B3))
M_i_5 net_0 B3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 VSS B2 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 net_0 B1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 ZN A1 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 net_0 A2 ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2 ZN A3 net_0 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_11 net_4 B3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_10 net_3 B2 net_4 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 ZN B1 net_3 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_1 A1 ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 net_2 A2 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 VDD A3 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR2_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:21:49 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR2_X1 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 + A2)
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_5 VDD A2 net_0 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR2_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:21:36 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR2_X2 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 + A2)
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5 VDD A2 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR2_X4.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:21:21 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR2_X4 A1 A2 ZN VDD VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VSS:G 
*.EQN ZN=(A1 + A2)
M_i_3__m0_x2__m1 ZN_neg A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0_x2__m1 VSS A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0_x2__m0 ZN_neg A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0_x2__m0 VSS A2 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_2 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_3 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m0_m2__m1 net_0__m0_0__m1 A2 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_m2__m1 ZN_neg A1 net_0__m0_0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_4__m0_m2__m0 net_0__m0_0__m0_0 A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0_m2__m0 VDD A2 net_0__m0_0__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_2 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR3_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:14:16 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR3_X1 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 + A2) + A3)
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_6 net_1 A2 net_0 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 VDD A3 net_1 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR3_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:14:13 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR3_X2 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 + A2) + A3)
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6 net_1 A2 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 VDD A3 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR3_X4.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:14:20 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR3_X4 A1 A2 A3 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VSS:G 
*.EQN ZN=((A1 + A2) + A3)
M_i_4__m0 ZN_neg A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 VSS A2 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 ZN_neg A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 VSS A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 ZN_neg A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m1 VSS A3 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7__m0 net_1__m0_0 A3 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_5__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 VDD A3 net_1__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR4_X1.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:08:17 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=(((A1 + A2) + A3) + A4)
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_7 net_1 A2 net_0 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_8 net_2 A3 net_1 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_9 VDD A4 net_2 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR4_X2.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:08:10 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR4_X2 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=(((A1 + A2) + A3) + A4)
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7 net_1 A2 net_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8 net_2 A3 net_1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9 VDD A4 net_2 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR4_X4.                                                          *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:08:21 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT OR4_X4 A1 A2 A3 A4 ZN VDD VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VSS:G 
*.EQN ZN=(((A1 + A2) + A3) + A4)
M_i_5__m0 ZN_neg A4 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m0 VSS A3 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m0 ZN_neg A2 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m0 VSS A1 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_2__m1 ZN_neg A1 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_3__m1 VSS A2 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_4__m1 ZN_neg A3 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5__m1 VSS A4 ZN_neg VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_9__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_6__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_7__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_8__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_9__m1 VDD A4 net_2__m1 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRS_X1.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:58:05 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRS_X1 D RN SE SI SN CK Q QN VDD VSS 
*.PININFO D:I RN:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_132 Q net_019 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_125 VSS net_017 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_119 net_019 net_017 net_018 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_114 net_018 RN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_101 net_016 SN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_106 net_017 net_013 net_016 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_28 VSS CK net_004 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_95 VSS RN net_015 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_77 net_012 net_007 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_71 VSS net_007 net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_66 net_011 RN net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_35 net_005 net_004 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_60 VSS SN net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_41 net_006 net_002 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 SI VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_12 net_002 SE net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_22 VSS D net_003 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_0 VSS SE net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_290 Q net_019 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_277 VDD net_017 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_284 VDD net_017 net_019 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_270 net_019 RN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_255 net_017 SN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_262 VDD net_013 net_017 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_165 VDD CK net_004 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_248 VDD RN net_026 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_234 net_026 net_017 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_228 VDD net_007 net_025 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_217 VDD net_007 net_010 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_211 net_010 RN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_172 net_005 net_004 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_203 VDD SN net_023 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_189 net_023 net_010 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_183 VDD net_002 net_022 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_159 VDD SI net_021 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_149 net_002 SE net_020 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_145 net_020 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_138 VDD SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRS_X2.                                                       *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:58:01 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRS_X2 D RN SE SI SN CK Q QN VDD VSS 
*.PININFO D:I RN:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_132_2 Q net_019 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_132 Q net_019 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_125 VSS net_017 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_125_68 VSS net_017 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_114 net_018 net_017 VSS VSS NMOS_VTL W=0.310000U L=0.050000U
M_i_119 net_019 RN net_018 VSS NMOS_VTL W=0.310000U L=0.050000U
M_i_106 net_017 SN net_016 VSS NMOS_VTL W=0.310000U L=0.050000U
M_i_101 net_016 net_013 VSS VSS NMOS_VTL W=0.310000U L=0.050000U
M_i_28 VSS CK net_004 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_95 VSS RN net_015 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_77 net_012 net_007 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_71 VSS net_007 net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_66 net_011 RN net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_35 net_005 net_004 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_60 VSS SN net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_41 net_006 net_002 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 SI VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_12 net_002 SE net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_22 VSS D net_003 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_0 VSS SE net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_290_11 Q net_019 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_290 Q net_019 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_277 VDD net_017 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_277_67 VDD net_017 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_284 VDD net_017 net_019 VDD PMOS_VTL W=0.485000U L=0.050000U
M_i_270 net_019 RN VDD VDD PMOS_VTL W=0.485000U L=0.050000U
M_i_255 net_017 SN VDD VDD PMOS_VTL W=0.485000U L=0.050000U
M_i_262 VDD net_013 net_017 VDD PMOS_VTL W=0.485000U L=0.050000U
M_i_165 VDD CK net_004 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_248 VDD RN net_026 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_234 net_026 net_017 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_228 VDD net_007 net_025 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_217 VDD net_007 net_010 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_211 net_010 RN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_172 net_005 net_004 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_203 VDD SN net_023 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_189 net_023 net_010 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_183 VDD net_002 net_022 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_159 VDD SI net_021 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_149 net_002 SE net_020 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_145 net_020 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_138 VDD SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFR_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:57:35 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFFR_X1 D RN SE SI CK Q QN VDD VSS 
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_0 VSS net_000 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_13 VSS net_003 net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_21 net_001 RN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_39 VSS net_009 net_004 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_83 net_011 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 net_005 net_011 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_62 net_008 net_006 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_77 VSS net_013 net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_56 VSS RN net_007 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_104 VSS SI net_014 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_100 net_014 SE net_013 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_89 net_012 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_110 net_015 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_116 VDD net_000 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_123 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_129 VDD net_003 net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_136 net_017 RN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_151 VDD net_000 net_017 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_157 net_018 net_009 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_209 net_011 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_167 VDD net_011 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_188 net_019 net_006 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_203 VDD net_013 net_020 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_174 net_006 net_009 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_181 VDD RN net_006 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_215 net_021 SI VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_226 net_022 SE net_013 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_230 VDD D net_022 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_236 net_015 SE VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFR_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:56:45 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFFR_X2 D RN SE SI CK Q QN VDD VSS 
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_13 VSS net_003 net_000 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7_145 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 Q net_003 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 VSS net_000 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_10 VSS net_000 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_21 net_001 RN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_39 VSS net_009 net_004 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_83 net_011 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 net_005 net_011 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_62 net_008 net_006 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_77 VSS net_013 net_010 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_56 VSS RN net_007 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_104 VSS SI net_014 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_100 net_014 SE net_013 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_89 net_012 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_110 net_015 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_129 VDD net_003 net_000 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_123_146 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_123 Q net_003 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_116 VDD net_000 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_116_1 VDD net_000 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_136 net_017 RN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_151 VDD net_000 net_017 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_157 net_018 net_009 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_209 net_011 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_167 VDD net_011 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_188 net_019 net_006 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_203 VDD net_013 net_020 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_174 net_006 net_009 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_181 VDD RN net_006 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_215 net_021 SI VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_226 net_022 SE net_013 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_230 VDD D net_022 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_236 net_015 SE VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFS_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:56:36 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFFS_X1 D SE SI SN CK Q QN VDD VSS 
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_0 VSS SE net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_21 VSS D net_003 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_11 net_002 SE net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 SI VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_27 VSS CK net_004 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_34 net_005 net_004 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_006 net_002 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_60 VSS SN net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_66 net_010 net_007 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_73 net_011 net_007 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_87 VSS net_015 net_013 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_93 net_014 SN VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_97 net_015 net_012 net_014 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_110 Q net_012 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_103 VSS net_015 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_116 VDD SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_123 net_016 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_127 net_002 SE net_016 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_137 VDD SI net_017 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_143 VDD CK net_004 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_150 net_005 net_004 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_157 net_018 net_002 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_172 VDD net_010 net_019 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_178 net_019 SN VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_189 VDD net_007 net_010 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_197 net_021 net_007 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_212 VDD net_015 net_022 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_218 net_015 SN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_224 VDD net_012 net_015 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_237 Q net_012 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_230 VDD net_015 QN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFS_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:56:22 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFFS_X2 D SE SI SN CK Q QN VDD VSS 
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_0 VSS SE net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_21 VSS D net_003 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_11 net_002 SE net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 SI VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_27 VSS CK net_004 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_34 net_005 net_004 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_006 net_002 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_60 VSS SN net_009 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_73 net_011 net_007 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_87 VSS net_015 net_013 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_66 net_010 net_007 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_93 net_014 SN net_015 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_97 VSS net_012 net_014 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_110_2 Q net_012 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_110 Q net_012 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_103 VSS net_015 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_103_26 VSS net_015 QN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_116 VDD SE net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_123 net_016 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_127 net_002 SE net_016 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_137 VDD SI net_017 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_143 VDD CK net_004 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_150 net_005 net_004 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_157 net_018 net_002 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_172 VDD net_010 net_019 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_178 net_019 SN VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_197 net_021 net_007 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_212 VDD net_015 net_022 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_189 VDD net_007 net_010 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_218 net_015 SN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_224 VDD net_012 net_015 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_237_1 Q net_012 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_237 Q net_012 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_230 VDD net_015 QN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_230_17 VDD net_015 QN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFF_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:55:24 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFF_X1 D SE SI CK Q QN VDD VSS 
*.PININFO D:I SE:I SI:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_7 QN net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 VSS net_002 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_13 VSS net_002 net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_20 net_001 net_000 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_34 VSS net_007 net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_004 net_009 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_75 net_009 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_54 net_006 net_005 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_69 VSS net_011 net_008 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_47 VSS net_007 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_96 VSS SI net_012 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_92 net_012 SE net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_81 net_010 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_102 net_013 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_115 QN net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_108 VDD net_002 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_121 VDD net_002 net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_128 net_014 net_000 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_143 VDD net_007 net_015 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_149 net_004 net_009 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_182 net_009 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_162 net_016 net_005 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_176 VDD net_011 net_017 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_155 VDD net_007 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_189 net_018 SI VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_200 net_019 SE net_011 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_204 VDD D net_019 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_210 net_013 SE VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFF_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:55:29 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT SDFF_X2 D SE SI CK Q QN VDD VSS 
*.PININFO D:I SE:I SI:I CK:I Q:O QN:O VDD:P VSS:G 
M_i_13 VSS net_002 net_000 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_50 VSS net_002 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 VSS net_002 Q VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 QN net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7_4 QN net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_20 net_001 net_000 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_34 VSS net_007 net_003 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_40 net_004 net_009 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_75 net_009 CK VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_54 net_006 net_005 VSS VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_69 VSS net_011 net_008 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_47 VSS net_007 net_005 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_96 VSS SI net_012 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_92 net_012 SE net_011 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_81 net_010 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_102 net_013 SE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_121 VDD net_002 net_000 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_108_51 VDD net_002 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_108 VDD net_002 Q VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_115 QN net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_115_2 QN net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_128 net_014 net_000 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_143 VDD net_007 net_015 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_149 net_004 net_009 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_182 net_009 CK VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_162 net_016 net_005 VDD VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_176 VDD net_011 net_017 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_155 VDD net_007 net_005 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_189 net_018 SI VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_200 net_019 SE net_011 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_204 VDD D net_019 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_210 net_013 SE VDD VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TBUF_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:21:14 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT TBUF_X1 A EN Z VDD VSS 
*.PININFO A:I EN:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_0 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_15_63 dummy1 A y VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0_15 VSS A x VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_0_14 VSS EN x VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_17 VSS EN NEN VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_24 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_0_64 VDD A y VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_24_1_48 y NEN VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_24_0 VDD A dummy0 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_24_1 dummy0 EN x VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_42 VDD EN NEN VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TBUF_X16.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:20:34 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT TBUF_X16 A EN Z VDD VSS 
*.PININFO A:I EN:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_0_6_6_40_125 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_13_45_122 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_37_112 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_42_108 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_6_43 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_13_120 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_106 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_116 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_13_45 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_37 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_42 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_6 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_13 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_63 dummy1a A y VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14_113 VSS EN x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_129 VSS A x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS A x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14 VSS EN x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17 VSS EN NEN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_24_3_19_50_12 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_8_39_66 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_18_103 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_9_17 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_19_51 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_8_42 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_83 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_10 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_8_39 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_18 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_9 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_19 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_8 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_1_48 y NEN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_64 VDD A y VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_64_92 VDD A y VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_130 x A dummy0a VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0 x A dummy0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_42 VDD EN NEN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TBUF_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:21:00 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT TBUF_X2 A EN Z VDD VSS 
*.PININFO A:I EN:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_0_6 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_14 VSS EN x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS A x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_63 dummy1 A y VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17 VSS EN NEN VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_24_3 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_1 dummy0 EN x VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0 VDD A dummy0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_64 VDD A y VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1_48 y NEN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_42 VDD EN NEN VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TBUF_X4.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:20:21 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT TBUF_X4 A EN Z VDD VSS 
*.PININFO A:I EN:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_0_6_6 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_13 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_63 dummy1 A y VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS A x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14 VSS EN x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17 VSS EN NEN VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_24_3_19 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_8 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_1_48 y NEN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_64 VDD A y VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0 x A dummy0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_42 VDD EN NEN VDD PMOS_VTL W=0.315000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TBUF_X8.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:20:37 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT TBUF_X8 A EN Z VDD VSS 
*.PININFO A:I EN:I Z:O VDD:P VSS:G 
*.EQN Z=A
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_13_45 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_37 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_42 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6_6 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_13 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_6 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0 VSS x Z VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_63 dummy1a A y VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14_113 VSS EN x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15_129 VSS A x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_15 VSS A x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0_14 VSS EN x VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17 VSS EN NEN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_8_39 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_18 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_9 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3_19 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_8 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_3 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24 VDD y Z VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_24_1_48 y NEN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_64 VDD A y VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_64_92 VDD A y VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0_130 x A dummy0a VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_0 x A dummy0 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_42 VDD EN NEN VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TINV_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:19:40 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT TINV_X1 EN I ZN VDD VSS 
*.PININFO EN:I I:I ZN:O VDD:P VSS:G 
*.EQN ZN=!I
M_i_0 VSS EN net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 I VSS VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_11 ZN net_000 net_001 VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_17 VDD EN net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_24 net_002 I VDD VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_29 ZN EN net_002 VDD PMOS_VTL W=0.540000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TLAT_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 18:55:08 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT TLAT_X1 D G OE Q VDD VSS 
*.PININFO D:I G:I OE:I Q:O VDD:P VSS:G 
M_i_0 VSS G net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 net_001 net_000 VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 net_002 D VSS VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL W=0.275000U L=0.050000U
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_28 VSS net_006 net_004 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_40 VSS net_003 net_006 VSS NMOS_VTL W=0.090000U L=0.050000U
M_i_34 net_005 OE VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_47 net_007 net_003 VSS VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_51 Q OE net_007 VSS NMOS_VTL W=0.355000U L=0.050000U
M_i_57 VDD G net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_64 net_001 net_000 VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_70 net_008 D VDD VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_75 net_003 net_000 net_008 VDD PMOS_VTL W=0.420000U L=0.050000U
M_i_81 net_009 net_001 net_003 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_85 VDD net_006 net_009 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_99 VDD net_003 net_006 VDD PMOS_VTL W=0.090000U L=0.050000U
M_i_91 net_005 OE VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_106 net_010 net_003 VDD VDD PMOS_VTL W=0.540000U L=0.050000U
M_i_111 Q net_005 net_010 VDD PMOS_VTL W=0.540000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR2_X1.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:19:40 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT XNOR2_X1 A B ZN VDD VSS 
*.PININFO A:I B:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A ^ B)
M_i_0 net_001 A net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_5 VSS B net_001 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_11 net_002 net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17 ZN A net_002 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_23 net_002 B ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_29 net_000 A VDD VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_36 VDD B net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_42 ZN net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_48 net_003 A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53 VDD B net_003 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR2_X2.                                                        *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:19:17 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT XNOR2_X2 A B ZN VDD VSS 
*.PININFO A:I B:I ZN:O VDD:P VSS:G 
*.EQN ZN=!(A ^ B)
M_i_11_23 net_002 net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_11 net_002 net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_5 VSS B net_001 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_0 net_001 A net_000 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17_20 ZN A net_002 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_17 ZN A net_002 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_23_12 net_002 B ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_23 net_002 B ZN VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_42_14 ZN net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_42 ZN net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_36 VDD B net_000 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_29 net_000 A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_48 net_003 A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_48_8 net_003b A ZN VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53_25 VDD B net_003b VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53 VDD B net_003 VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR2_X1.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:19:03 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT XOR2_X1 A B Z VDD VSS 
*.PININFO A:I B:I Z:O VDD:P VSS:G 
*.EQN Z=(A ^ B)
M_i_0 net_000 A VSS VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_7 VSS B net_000 VSS NMOS_VTL W=0.210000U L=0.050000U
M_i_13 Z net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_19 net_001 A Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_24 VSS B net_001 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_30 net_002 A net_000 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_35 VDD B net_002 VDD PMOS_VTL W=0.315000U L=0.050000U
M_i_41 net_003 net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_47 Z A net_003 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53 net_003 B Z VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR2_X2.                                                         *
*                                                                              *
* Technology: NCSU FreePDK 45nm.                                               *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr)     *
* at 19:19:07 on Fri, 3 Dec 2010.                                              *
*                                                                              *
********************************************************************************
.SUBCKT XOR2_X2 A B Z VDD VSS 
*.PININFO A:I B:I Z:O VDD:P VSS:G 
*.EQN Z=(A ^ B)
M_i_0 net_000 A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_7 VSS B net_000 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_13 Z net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_19 net_001 A Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_24 VSS B net_001 VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_24_4 VSS B net_001b VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_19_23 net_001b A Z VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_13_35 Z net_000 VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_30 net_002 A net_000 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_35 VDD B net_002 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_41 net_003 net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_47 Z A net_003 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53 net_003 B Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_53_18 net_003 B Z VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_47_27 Z A net_003 VDD PMOS_VTL W=0.630000U L=0.050000U
M_i_41_29 net_003 net_000 VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
